----------------------------------------------------------------------------------
-- Company: UFSJ
-- Engineer: Nathan Lima
-- 
-- Create Date:    07:59:36 01/24/2025 
-- Design Name: 
-- Module Name:    deslocador_2b_esq - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity deslocador_2b_esq is
    port(
        entrada: in std_logic_vector(31 downto 0);
        saida: out std_logic_vector(31 downto 0)
    );
end deslocador_2b_esq;

architecture Behavioral of deslocador_2b_esq is
begin
    process(entrada)
    begin
        saida(31 downto 2) <= entrada(29 downto 0);
        saida(1 downto 0) <= "00";
    end process;
end Behavioral;
